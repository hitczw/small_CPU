module CPU_top(RST,CLK,ACCUM_OUT);
input RST;
input CLK;

wire[7:0] DATA;
wire[2:0] OPCODE;
wire[12:0] IR_ADDR;
wire LOAD_IR;

output wire[7:0] ACCUM_OUT;


wire[7:0] ACCUM_IN;
wire LOAD_ACC;

wire ZERO;

wire FETCH;
wire INC_PC;
wire LOAD_PC;
wire RD;
wire WR;
wire DATACTL_ENA;

wire[12:0] PC_ADDR;
wire[12:0] ADDR;

wire ALU_N;
wire ALU_ENA;
wire[7:0] ALU_OUT;


//REGISTER(DATA,ENA,CLK,OPCODE,IR_ADDR);
REGISTER re(DATA,LOAD_IR,CLK,OPCODE,IR_ADDR);

//ACCUMULATOR(ALU_OUT,LOAD_ACC,RST,ACCUM,ZERO);
ACCUMULATOR ac(ACCUM_IN,LOAD_ACC,RST,ACCUM_OUT,ZERO);

//ALU(DATA,ACCUM,OPCODE,ALU_OUT);
ALU al(DATA,ACCUM_OUT,OPCODE,ALU_OUT,ALU_ENA,CLK);

//module CONTROL(CLK1,RST,OPCODE,ZERO,INC_PC,LOAD_ACC,LOAD_PC,RD,WD,LOAD_IR,DATACTL_ENA,ALU_CLOCK,FETCH,ALU_N);
CONTROL co(CLK,RST,OPCODE,ZERO,INC_PC,LOAD_ACC,LOAD_PC,RD,WR,LOAD_IR,DATACTL_ENA,FETCH,ALU_N,ALU_ENA);

//module DATACTL(IN,DATA_ENA,DATA);
DATACTL da(ACCUM_OUT,DATACTL_ENA,DATA);

//ADDR(FETCH,IR_ADDR,PC_ADDR,OUT_ADDR);
ADDR ad(FETCH,IR_ADDR,PC_ADDR,ADDR);

//COUNTER(IR_ADDR,LOAD,CLOCK,RST,OUT_ADDR);
COUNTER cou(IR_ADDR,LOAD_PC,INC_PC,RST,PC_ADDR);

//module CHOOSE(IR_ADDR,ALU_OUT,ALU_N,OUT_DATA);
CHOOSE ch(IR_ADDR,ALU_OUT,ALU_N,ACCUM_IN);

//RAOM(data,addr,read,write);
RAOM ra(DATA,ADDR,RD,WR);


endmodule